module	Lab1_gatelevel_UDP(F, A, B, C);
	output	F;
	input	A, B, C;

	Lab1_UDP M0(F, A, B, C);

endmodule